* SPICE NETLIST
***************************************

.SUBCKT mim_cap_test A B
** N=2 EP=2 IP=0 FDC=1
C0 A B area=4e-10 perimeter=8e-05 $[cmmh4] $X=-1245 $Y=-1245 $D=0
.ENDS
***************************************
