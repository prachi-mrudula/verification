* SPICE NETLIST
***************************************

.SUBCKT qpva5
** N=3 EP=0 IP=0 FDC=1
Q0 1 2 3 qpva5 $X=3150 $Y=3150 $D=0
.ENDS
***************************************
