* SPICE NETLIST
***************************************

.SUBCKT res_test A B
** N=155 EP=2 IP=0 FDC=1
R0 A B L=1e-05 W=2e-06 $[rnp1] $X=-1025 $Y=-1525 $D=0
.ENDS
***************************************
