* SPICE NETLIST
***************************************

.SUBCKT PE_5 D G S B SB
.ENDS
***************************************
.SUBCKT PEL_5 D G S B SB
.ENDS
***************************************
.SUBCKT PESVT_5 D G S B SB
.ENDS
***************************************
.SUBCKT MOSVC G NW SB
.ENDS
***************************************
.SUBCKT MOSVCTI G PW
.ENDS
***************************************
.SUBCKT LDDN D G S B
.ENDS
***************************************
.SUBCKT LDDP D G S B
.ENDS
***************************************
.SUBCKT MOSVC5 G NW SB
.ENDS
***************************************
.SUBCKT MOSVC5TI G PW
.ENDS
***************************************
.SUBCKT NHSJ1_7 D G S B HW
.ENDS
***************************************
.SUBCKT NHSJ1_10 D G S B HW
.ENDS
***************************************
.SUBCKT NHSJ1_16C D G S B HW
.ENDS
***************************************
.SUBCKT PHSJ1_7 D G S B HW
.ENDS
***************************************
.SUBCKT PHSJ1_10 D G S B HW
.ENDS
***************************************
.SUBCKT PHSJ1_16C D G S B HW
.ENDS
***************************************
.SUBCKT PE5_5 D G S B SB
.ENDS
***************************************
.SUBCKT NHVTA D G S B HW
.ENDS
***************************************
.SUBCKT NHVTAA D G S B HW
.ENDS
***************************************
.SUBCKT NHVTB D G S B HW
.ENDS
***************************************
.SUBCKT NHVU D G S B HW
.ENDS
***************************************
.SUBCKT NDHVT D G S B HW
.ENDS
***************************************
.SUBCKT NDHVTA D G S B HW
.ENDS
***************************************
.SUBCKT NDHVTAA D G S B HW
.ENDS
***************************************
.SUBCKT PHVTA D G S B HW
.ENDS
***************************************
.SUBCKT PHVTB D G S B HW
.ENDS
***************************************
.SUBCKT PHVU D G S B HW
.ENDS
***************************************
.SUBCKT NMVB D G S B HW
.ENDS
***************************************
.SUBCKT NMVC D G S B HW
.ENDS
***************************************
.SUBCKT NMVD D G S B HW
.ENDS
***************************************
.SUBCKT NMVE D G S B HW
.ENDS
***************************************
.SUBCKT NMVF D G S B HW
.ENDS
***************************************
.SUBCKT NDMVD D G S B HW
.ENDS
***************************************
.SUBCKT NDMVF D G S B HW
.ENDS
***************************************
.SUBCKT PMVB D G S B HW
.ENDS
***************************************
.SUBCKT PMVC D G S B HW
.ENDS
***************************************
.SUBCKT PMVD D G S B HW
.ENDS
***************************************
.SUBCKT PMVE D G S B HW
.ENDS
***************************************
.SUBCKT PMVF D G S B HW
.ENDS
***************************************
.SUBCKT NHVRA D G S B HW
.ENDS
***************************************
.SUBCKT NHVRB D G S B HW
.ENDS
***************************************
.SUBCKT NHVRC D G S B HW
.ENDS
***************************************
.SUBCKT NHVRD D G S B HW
.ENDS
***************************************
.SUBCKT NHVRE D G S B HW
.ENDS
***************************************
.SUBCKT NHVRF D G S B HW
.ENDS
***************************************
.SUBCKT NDHVRD D G S B HW
.ENDS
***************************************
.SUBCKT NDHVRF D G S B HW
.ENDS
***************************************
.SUBCKT PHVRA D G S B HW
.ENDS
***************************************
.SUBCKT PHVRB D G S B HW
.ENDS
***************************************
.SUBCKT PHVRC D G S B HW
.ENDS
***************************************
.SUBCKT PHVRD D G S B HW
.ENDS
***************************************
.SUBCKT PHVRE D G S B HW
.ENDS
***************************************
.SUBCKT PHVRF D G S B HW
.ENDS
***************************************
.SUBCKT NISJ1_16 C G E HW
.ENDS
***************************************
.SUBCKT tag_200v N1
.ENDS
***************************************
.SUBCKT tag_100v N1
.ENDS
***************************************
.SUBCKT tag_60v N1
.ENDS
***************************************
.SUBCKT tag_25v N1
.ENDS
***************************************
.SUBCKT tag_m200v N1
.ENDS
***************************************
.SUBCKT tag_m100v N1
.ENDS
***************************************
.SUBCKT tag_m60v N1
.ENDS
***************************************
.SUBCKT tag_m25v N1
.ENDS
***************************************
.SUBCKT ne5_m2 G B D S
** N=5 EP=4 IP=0 FDC=2
M0 S G D B ne5 L=5e-07 W=2e-06 AD=5.4e-13 AS=9.6e-13 PD=2.54e-06 PS=4.96e-06 $X=27195 $Y=-1380 $D=13
M1 D G S B ne5 L=5e-07 W=2e-06 AD=9.6e-13 AS=5.4e-13 PD=4.96e-06 PS=2.54e-06 $X=28235 $Y=-1380 $D=13
.ENDS
***************************************
