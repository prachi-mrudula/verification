* SPICE NETLIST
***************************************

.SUBCKT pe_test B G S D
** N=97 EP=4 IP=0 FDC=1
M0 D G S B pe L=1.8e-07 W=2e-06 AD=9.6e-13 AS=9.6e-13 PD=4.96e-06 PS=4.96e-06 $X=8350 $Y=-4375 $D=0
.ENDS
***************************************
