* SPICE NETLIST
***************************************

.SUBCKT res_create
** N=82 EP=0 IP=0 FDC=1
R0 38 22 L=1.70505e-06 W=6.0825e-06 $[rnp1] $X=11080 $Y=10855 $D=0
.ENDS
***************************************
