* SPICE NETLIST
***************************************

.SUBCKT rnw_test C A B
** N=3 EP=3 IP=0 FDC=1
R0 A B L=1e-05 W=2e-06 $SUB=C $[rnw5] $X=-605 $Y=-1145 $D=0
.ENDS
***************************************
