* SPICE NETLIST
***************************************

.SUBCKT ser_res_test1 A B C D
** N=4 EP=4 IP=0 FDC=2
R0 A B L=0.00387656 W=2e-05 $[rnp1] $X=-1025 $Y=-1525 $D=0
R1 C D L=0.00387656 W=2e-05 $[rnp1] $X=524385 $Y=322665 $D=0
.ENDS
***************************************
