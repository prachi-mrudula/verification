* SPICE NETLIST
***************************************

.SUBCKT ser_res_test A B
** N=403 EP=2 IP=0 FDC=1
R0 A B L=0.00030762 W=2e-06 $[rnp1] $X=-1025 $Y=-1525 $D=0
.ENDS
***************************************
