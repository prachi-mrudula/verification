* SPICE NETLIST
***************************************

.SUBCKT ser_45_test C D
** N=2 EP=2 IP=0 FDC=1
R0 C D L=6.11674e-05 W=2e-06 $[rnp1] $X=-1025 $Y=-1525 $D=0
.ENDS
***************************************
